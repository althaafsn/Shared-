







task automatic taskName();
    
endtask //automatic

