module cpuTest();

    







endmodule