

module regfile_tb();
    
endmodule